`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 09/12/2023 03:55:15 PM
// Design Name: 
// Module Name: AXI_top_tb
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// Based on: https://www.realdigital.org/doc/32101c99686fe25ec47bedd94e76dc96
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module AXI_top_tb();
//clock and reset_n signals

    parameter reg0_addr = 32'b0;
    parameter reg1_addr = 32'h00000004;
	parameter reg2_addr = 32'h00000008;
	parameter reg3_addr = 32'h0000000c;
    
    
    
    
	reg aclk =1'b0;
	reg arstn = 1'b0;

	
	//Write Address channel (AW)
	reg [31:0] write_addr =32'd0;	//Master write address
	reg [2:0] write_prot = 3'd0;	//type of write(leave at 0)
	reg write_addr_valid = 1'b0;	//master indicating address is valid
	wire write_addr_ready;		//slave ready to receive address

	//Write Data Channel (W)
	reg [31:0] write_data = 32'd0;	//Master write data
	reg [3:0] write_strb = 4'd0;	//Master byte-wise write strobe
	reg write_data_valid = 1'b0;	//Master indicating write data is valid
	wire write_data_ready;		//slave ready to receive data

	//Write Response Channel (WR)
	reg write_resp_ready = 1'b0;	//Master ready to receive write response
	wire [1:0] write_resp;		//slave write response
	wire write_resp_valid;		//slave response valid
	
	//Read Address channel (AR)
	reg [31:0] read_addr = 32'd0;	//Master read address
	reg [2:0] read_prot =3'd0;	//type of read(leave at 0)
	reg read_addr_valid = 1'b0;	//Master indicating address is valid
	wire read_addr_ready;		//slave ready to receive address

	//Read Data Channel (R)
	reg read_data_ready = 1'b0;	//Master indicating ready to receive data
	wire [31:0] read_data;		//slave read data
	wire [1:0] read_resp;		//slave read response
	wire read_data_valid;		//slave indicating data in channel is valid 
    
    BCP_accelerator_v2_0_S01_AXI #(
        .C_S_AXI_DATA_WIDTH(32),
		.C_S_AXI_ADDR_WIDTH(32)
    )DUT(
		.S_AXI_ACLK(aclk),
		.S_AXI_ARESETN(arstn),

		.S_AXI_AWADDR(write_addr),
		.S_AXI_AWPROT(write_prot),
		.S_AXI_AWVALID(write_addr_valid),
		.S_AXI_AWREADY(write_addr_ready),

		.S_AXI_WDATA(write_data),
		.S_AXI_WSTRB(write_strb),
		.S_AXI_WVALID(write_data_valid),
		.S_AXI_WREADY(write_data_ready),

		.S_AXI_BRESP(write_resp),
		.S_AXI_BVALID(write_resp_valid),
		.S_AXI_BREADY(write_resp_ready),

		.S_AXI_ARADDR(read_addr),
		.S_AXI_ARPROT(read_prot),
		.S_AXI_ARVALID(read_addr_valid),
		.S_AXI_ARREADY(read_addr_ready),

		.S_AXI_RDATA(read_data),
		.S_AXI_RRESP(read_resp),
		.S_AXI_RVALID(read_data_valid),
		.S_AXI_RREADY(read_data_ready)
    );
    
    always 
        #5 aclk <= ~aclk;
        
    integer i;	
	initial
	begin
   		arstn = 0;
		i=0;
		#20 arstn=1;
		
		// Write clause to FPGA
		//		for(i=0;i<=32'hF;i=i+1)	
        //      #20 axi_write(32'd0,i);	//write i to slv_reg0\
		update_clause(30'd0,32'd8,1'b1,32'd9,1'b0,32'd7,1'b1); // 8 -9 7 SAT
		#60;
        update_clause(30'd1,32'd7,1'b0,32'd9,1'b1,32'd15,1'b0); // -7 9 -15 SAT
		#60;
		update_clause(30'd2,32'd9,1'b1,32'd8,1'b1,32'd1,1'b1); // 9 8 1 SAT
		#60;
		update_clause(30'd3,32'd5,1'b1,32'd19,1'b1,32'd2,1'b1); // 5 -19 2 
		#60;
		update_clause(30'd4,32'd1,1'b0,32'd9,1'b0,32'd8,1'b0); // -1 -9 -8 SAT
		#60;
		update_clause(30'd5,32'd4,1'b1,32'd19,1'b1,32'd16,1'b1); // 4 19 16
		#60;
		
		// Send Decision to FPGA
		send_decision(1'b0,30'd1,1'b0); // No changes to status, Clause 4 is now SAT
		send_decision(1'b0,30'd9,1'b0); // Unit implication generated by clause 2 (var id 8, polarity = 1), Clause 0 now SAT, Clause 2 now SAT
		
		// Backtrack and remove unit implication (this should never happen, but I want to test the system running into a conflict state)
		send_decision(1'b1,30'd8,1'b0);
//		send_decision(1'b1,30'd9,1'b0); // Unit implication generated by clause 2 (var id 8, polarity = 1), Clause 0 now SAT, Clause 2 now SAT
		// Create conflict
		send_decision(1'b0,30'd8,1'b0);
		send_decision(1'b1,30'd8,1'b0);
		
		// Create SAT
		send_decision(1'b0,30'd9,1'b0); // 0, 4 and 2 now SAT
		send_decision(1'b0,30'd7,1'b0); // 1 now SAT
		send_decision(1'b0,30'd2,1'b1); // 3 now SAT
		send_decision(1'b0,30'd19,1'b1); // 0, 4 and 2 now SAT
		
		
		#500;
		$finish;
	end
	
	task axi_write;
	input [31:0] addr;
	input [31:0] data;
	begin
		#3 write_addr <= addr;	//Put write address on bus
		write_data <= data;	//put write data on bus
		write_addr_valid <= 1'b1;	//indicate address is valid
		write_data_valid <= 1'b1;	//indicate data is valid
		write_resp_ready <= 1'b1;	//indicate ready for a response
		write_strb <= 4'hF;		//writing all 4 bytes

		//wait for one slave ready signal or the other
		wait(write_data_ready || write_addr_ready);
			
		@(posedge aclk); //one or both signals and a positive edge
		if(write_data_ready&&write_addr_ready)//received both ready signals
		begin
			write_addr_valid<=0;
			write_data_valid<=0;
		end
		else    //wait for the other signal and a positive edge
		begin
			if(write_data_ready)    //case data handshake completed
			begin
				write_data_valid<=0;
				wait(write_addr_ready); //wait for address address ready
			end
            		else if(write_addr_ready)   //case address handshake completed
            		begin
				write_addr_valid<=0;
                		wait(write_data_ready); //wait for data ready
            		end 
			@ (posedge aclk);// complete the second handshake
			write_addr_valid<=0; //make sure both valid signals are deasserted
			write_data_valid<=0;
		end
            
		//both handshakes have occured
		//deassert strobe
		write_strb<=0;

		//wait for valid response
		wait(write_resp_valid);
		
		//both handshake signals and rising edge
		@(posedge aclk);

		//deassert ready for response
		write_resp_ready<=0;

		//end of write transaction
	end
	endtask;
	
	task update_clause;
	input [29:0] clause_id;
	input [30:0] var1;
	input        var1_pol;
	input [30:0] var2;
	input        var2_pol;
	input [30:0] var3;
	input        var3_pol;
	begin
	   #20 axi_write(32'd0,32'h00000000);
	   // Write reg1;
	   #20 axi_write(32'h00000004,{var1,var1_pol});
	   // write reg2;
	   #20 axi_write(32'h00000008,{var2,var2_pol});
	   // write reg3;
	   #20 axi_write(32'h0000000c,{var3,var3_pol});
	   //write reg 0;
	   #20 axi_write(32'h0,{clause_id,2'b01}); // Update clause ID OP code = 001
	end;
	endtask;
	
	task send_decision;
	input backtrack;
	input [30:0] var_id;
	input        decision_polarity;
	begin
	   #20 axi_write(reg0_addr, 32'd0);
	   // Write reg 1
	   #20 axi_write(reg1_addr, {var_id,decision_polarity});
	   // Write reg 0 with CPU OP code 10
	   if(backtrack) begin
	       #20 axi_write(reg0_addr,32'h00000003);
	   end else begin
	       #20 axi_write(reg0_addr,32'h00000002);
	   end
	   // Verify
	end
	endtask

endmodule
